module moduleName (instrucao, saida);
    input [31:0] instrucao;
    output reg[31:0] saida;

    
endmodule