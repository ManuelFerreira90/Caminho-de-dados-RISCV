module memoria (clk, aluresult2, rs2, reddataM, memwrite, memread, immediate, mem0, mem1, mem2, mem3, mem4, mem5, mem6, mem7, mem8, mem9, mem10, mem11, mem12, mem13, mem14, mem15, mem16, mem17, mem18, mem19, mem20, mem21, mem22, mem23, mem24, mem25, mem26, mem27, mem28, mem29, mem30, mem31, mem32, mem33, mem34, mem35, mem36, mem37, mem38, mem39, mem40, mem41, mem42, mem43, mem44, mem45, mem46, mem47, mem48, mem49, mem50, mem51, mem52, mem53, mem54, mem55, mem56, mem57, mem58, mem59, mem60, mem61, mem62, mem63, estado);
    input wire clk;
    input [2:0] estado;   
    input [31:0] aluresult2;
    input [4:0] rs2;
    input memwrite;
    input memread;
    input [11:0] immediate;
    output reg [31:0] reddataM;
    output reg [31:0] mem0, mem1, mem2, mem3, mem4, mem5, mem6, mem7, mem8, mem9, mem10, mem11;
    output reg [31:0] mem12, mem13, mem14, mem15, mem16, mem17, mem18, mem19, mem20, mem21, mem22, mem23; 
    output reg [31:0] mem24, mem25, mem26, mem27, mem28, mem29, mem30, mem31, mem32, mem33, mem34, mem35, mem36, mem37, mem38, mem39, mem40, mem41, mem42, mem43, mem44, mem45, mem46, mem47, mem48, mem49, mem50, mem51, mem52, mem53, mem54, mem55, mem56, mem57, mem58, mem59, mem60, mem61, mem62, mem63;
    //reg [31:0] immediateaux;
    reg [63:0] memoria [0:63];

    initial begin
        $readmemb("entrada/memoria.bin", memoria); // iniciando a memoria
        mem0 <= memoria[0];
        mem1 <= memoria[1];
        mem2 <= memoria[2];
        mem3 <= memoria[3];
        mem4 <= memoria[4];
        mem5 <= memoria[5];
        mem6 <= memoria[6];
        mem7 <= memoria[7];
        mem8 <= memoria[8];
        mem9 <= memoria[9];
        mem10 <= memoria[10];
        mem11 <= memoria[11];
        mem12 <= memoria[12];
        mem13 <= memoria[13];
        mem14 <= memoria[14];
        mem15 <= memoria[15];
        mem16 <= memoria[16];
        mem17 <= memoria[17];
        mem18 <= memoria[18];
        mem19 <= memoria[19];
        mem20 <= memoria[20];
        mem21 <= memoria[21];
        mem22 <= memoria[22];
        mem23 <= memoria[23];
        mem24 <= memoria[24];
        mem25 <= memoria[25];
        mem26 <= memoria[26];
        mem27 <= memoria[27];
        mem28 <= memoria[28];
        mem29 <= memoria[29];
        mem30 <= memoria[30];
        mem31 <= memoria[31];
        mem32 <= memoria[32];  
        mem33 <= memoria[33];  
        mem34 <= memoria[34];  
        mem35 <= memoria[35];  
        mem36 <= memoria[36];  
        mem37 <= memoria[37];  
        mem38 <= memoria[38];  
        mem39 <= memoria[39];  
        mem40 <= memoria[40];  
        mem41 <= memoria[41];  
        mem42 <= memoria[42];  
        mem43 <= memoria[43];  
        mem44 <= memoria[44];  
        mem45 <= memoria[45];  
        mem46 <= memoria[46];  
        mem47 <= memoria[47];  
        mem48 <= memoria[48];  
        mem49 <= memoria[49];  
        mem50 <= memoria[50];  
        mem51 <= memoria[51];  
        mem52 <= memoria[52];  
        mem53 <= memoria[53];  
        mem54 <= memoria[54];  
        mem55 <= memoria[55];  
        mem56 <= memoria[56];  
        mem57 <= memoria[57];  
        mem58 <= memoria[58];  
        mem59 <= memoria[59];  
        mem60 <= memoria[60];  
        mem61 <= memoria[61];  
        mem62 <= memoria[62];   
        mem63 <= memoria[63];
    end

    always @(posedge clk) begin
        //immediateaux <= immediate / 4;
        if(estado == 3'b100) begin
            if(memwrite == 1'b1) begin
                memoria[aluresult2] <= rs2;
            end
            if(memread == 1'b1) begin
                reddataM <= memoria[aluresult2];
            end
            mem0 <= memoria[0];
            mem1 <= memoria[1];
            mem2 <= memoria[2];
            mem3 <= memoria[3];
            mem4 <= memoria[4];
            mem5 <= memoria[5];
            mem6 <= memoria[6];
            mem7 <= memoria[7];
            mem8 <= memoria[8];
            mem9 <= memoria[9];
            mem10 <= memoria[10];
            mem11 <= memoria[11];
            mem12 <= memoria[12];
            mem13 <= memoria[13];
            mem14 <= memoria[14];
            mem15 <= memoria[15];
            mem16 <= memoria[16];
            mem17 <= memoria[17];
            mem18 <= memoria[18];
            mem19 <= memoria[19];
            mem20 <= memoria[20];
            mem21 <= memoria[21];
            mem22 <= memoria[22];
            mem23 <= memoria[23];
            mem24 <= memoria[24];
            mem25 <= memoria[25];
            mem26 <= memoria[26];
            mem27 <= memoria[27];
            mem28 <= memoria[28];
            mem29 <= memoria[29];
            mem30 <= memoria[30];
            mem31 <= memoria[31];     
            mem32 <= memoria[32];  
            mem33 <= memoria[33];  
            mem34 <= memoria[34];  
            mem35 <= memoria[35];  
            mem36 <= memoria[36];  
            mem37 <= memoria[37];  
            mem38 <= memoria[38];  
            mem39 <= memoria[39];  
            mem40 <= memoria[40];  
            mem41 <= memoria[41];  
            mem42 <= memoria[42];  
            mem43 <= memoria[43];  
            mem44 <= memoria[44];  
            mem45 <= memoria[45];  
            mem46 <= memoria[46];  
            mem47 <= memoria[47];  
            mem48 <= memoria[48];  
            mem49 <= memoria[49];  
            mem50 <= memoria[50];  
            mem51 <= memoria[51];  
            mem52 <= memoria[52];  
            mem53 <= memoria[53];  
            mem54 <= memoria[54];  
            mem55 <= memoria[55];  
            mem56 <= memoria[56];  
            mem57 <= memoria[57];  
            mem58 <= memoria[58];  
            mem59 <= memoria[59];  
            mem60 <= memoria[60];  
            mem61 <= memoria[61];  
            mem62 <= memoria[62];   
            mem63 <= memoria[63];  
        end
    end
    
endmodule