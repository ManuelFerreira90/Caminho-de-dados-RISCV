module alusrc (immediate, rs2);
    input wire immediate;
    
endmodule