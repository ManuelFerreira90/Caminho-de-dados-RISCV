module lerinstrucao (instrucao, pc, clk, estado, rst);
    input wire [31:0] pc;
    input clk, rst;
    input wire [3:0] estado;
    output reg [31:0] instrucao;
    // alterar confome a quantidade de linhas do arquivo
    reg [31:0] instrucoes [0:15]; // Memória de instruções

    // Atualizando instrução a cada ciclo de clock
    always @(posedge clk) begin
        if(rst == 1'b1) begin
            instrucoes [0] <= 32'b00000000011100000000000100010011;
				instrucoes [1] <= 32'b00000000001000000010001000100011;
				instrucoes [2] <= 32'b00000000010000000010000010000011;
				instrucoes [3] <= 32'b00000000000000001000000100110011;
				instrucoes [4] <= 32'b00000000001000001000000010110011;
				instrucoes [5] <= 32'b00000000001000001000000010110011;
				instrucoes [6] <= 32'b01000000001000001000000010110011;
				instrucoes [7] <= 32'b01000000001000001000000010110011;
				instrucoes [8] <= 32'b00000000001000001000011001100011;
				instrucoes [9] <= 32'b00000000000100001000000010110011;
				instrucoes [10] <= 32'b00000000000100000010000000100011;
				instrucoes [11] <= 32'b00000000001000001111000010110011;
				instrucoes [12] <= 32'b00000000000000001110000010110011;
				instrucoes [13] <= 32'b00000000000100000010000000100011;
				instrucoes [14] <= 32'b00000000000000000000000000000000;
				instrucoes [15] <= 32'b00000000000000000000000000000000;
        end
        if(estado == 4'b0000)begin
            instrucao <= instrucoes[pc];
        end
    end

endmodule


